`ifndef LINEARIZE_SVH
`define LINEARIZE_SVH

function logic [7:0] linearize(input logic [7:0] rgb);
    unique case (rgb)
        8'd0:   linearize = 8'd0;
        8'd1:   linearize = 8'd0;
        8'd2:   linearize = 8'd0;
        8'd3:   linearize = 8'd0;
        8'd4:   linearize = 8'd0;
        8'd5:   linearize = 8'd0;
        8'd6:   linearize = 8'd0;
        8'd7:   linearize = 8'd0;
        8'd8:   linearize = 8'd0;
        8'd9:   linearize = 8'd0;
        8'd10:  linearize = 8'd0;
        8'd11:  linearize = 8'd0;
        8'd12:  linearize = 8'd0;
        8'd13:  linearize = 8'd0;
        8'd14:  linearize = 8'd0;
        8'd15:  linearize = 8'd0;
        8'd16:  linearize = 8'd0;
        8'd17:  linearize = 8'd0;
        8'd18:  linearize = 8'd0;
        8'd19:  linearize = 8'd0;
        8'd20:  linearize = 8'd0;
        8'd21:  linearize = 8'd0;
        8'd22:  linearize = 8'd0;
        8'd23:  linearize = 8'd0;
        8'd24:  linearize = 8'd0;
        8'd25:  linearize = 8'd0;
        8'd26:  linearize = 8'd0;
        8'd27:  linearize = 8'd0;
        8'd28:  linearize = 8'd1;
        8'd29:  linearize = 8'd1;
        8'd30:  linearize = 8'd1;
        8'd31:  linearize = 8'd1;
        8'd32:  linearize = 8'd1;
        8'd33:  linearize = 8'd1;
        8'd34:  linearize = 8'd1;
        8'd35:  linearize = 8'd1;
        8'd36:  linearize = 8'd1;
        8'd37:  linearize = 8'd1;
        8'd38:  linearize = 8'd1;
        8'd39:  linearize = 8'd1;
        8'd40:  linearize = 8'd1;
        8'd41:  linearize = 8'd2;
        8'd42:  linearize = 8'd2;
        8'd43:  linearize = 8'd2;
        8'd44:  linearize = 8'd2;
        8'd45:  linearize = 8'd2;
        8'd46:  linearize = 8'd2;
        8'd47:  linearize = 8'd2;
        8'd48:  linearize = 8'd2;
        8'd49:  linearize = 8'd3;
        8'd50:  linearize = 8'd3;
        8'd51:  linearize = 8'd3;
        8'd52:  linearize = 8'd3;
        8'd53:  linearize = 8'd3;
        8'd54:  linearize = 8'd3;
        8'd55:  linearize = 8'd3;
        8'd56:  linearize = 8'd4;
        8'd57:  linearize = 8'd4;
        8'd58:  linearize = 8'd4;
        8'd59:  linearize = 8'd4;
        8'd60:  linearize = 8'd4;
        8'd61:  linearize = 8'd5;
        8'd62:  linearize = 8'd5;
        8'd63:  linearize = 8'd5;
        8'd64:  linearize = 8'd5;
        8'd65:  linearize = 8'd6;
        8'd66:  linearize = 8'd6;
        8'd67:  linearize = 8'd6;
        8'd68:  linearize = 8'd6;
        8'd69:  linearize = 8'd7;
        8'd70:  linearize = 8'd7;
        8'd71:  linearize = 8'd7;
        8'd72:  linearize = 8'd7;
        8'd73:  linearize = 8'd8;
        8'd74:  linearize = 8'd8;
        8'd75:  linearize = 8'd8;
        8'd76:  linearize = 8'd9;
        8'd77:  linearize = 8'd9;
        8'd78:  linearize = 8'd9;
        8'd79:  linearize = 8'd10;
        8'd80:  linearize = 8'd10;
        8'd81:  linearize = 8'd10;
        8'd82:  linearize = 8'd11;
        8'd83:  linearize = 8'd11;
        8'd84:  linearize = 8'd11;
        8'd85:  linearize = 8'd12;
        8'd86:  linearize = 8'd12;
        8'd87:  linearize = 8'd13;
        8'd88:  linearize = 8'd13;
        8'd89:  linearize = 8'd13;
        8'd90:  linearize = 8'd14;
        8'd91:  linearize = 8'd14;
        8'd92:  linearize = 8'd15;
        8'd93:  linearize = 8'd15;
        8'd94:  linearize = 8'd16;
        8'd95:  linearize = 8'd16;
        8'd96:  linearize = 8'd17;
        8'd97:  linearize = 8'd17;
        8'd98:  linearize = 8'd18;
        8'd99:  linearize = 8'd18;
        8'd100: linearize = 8'd19;
        8'd101: linearize = 8'd19;
        8'd102: linearize = 8'd20;
        8'd103: linearize = 8'd20;
        8'd104: linearize = 8'd21;
        8'd105: linearize = 8'd21;
        8'd106: linearize = 8'd22;
        8'd107: linearize = 8'd22;
        8'd108: linearize = 8'd23;
        8'd109: linearize = 8'd24;
        8'd110: linearize = 8'd24;
        8'd111: linearize = 8'd25;
        8'd112: linearize = 8'd25;
        8'd113: linearize = 8'd26;
        8'd114: linearize = 8'd27;
        8'd115: linearize = 8'd27;
        8'd116: linearize = 8'd28;
        8'd117: linearize = 8'd29;
        8'd118: linearize = 8'd29;
        8'd119: linearize = 8'd30;
        8'd120: linearize = 8'd31;
        8'd121: linearize = 8'd32;
        8'd122: linearize = 8'd32;
        8'd123: linearize = 8'd33;
        8'd124: linearize = 8'd34;
        8'd125: linearize = 8'd35;
        8'd126: linearize = 8'd35;
        8'd127: linearize = 8'd36;
        8'd128: linearize = 8'd37;
        8'd129: linearize = 8'd38;
        8'd130: linearize = 8'd39;
        8'd131: linearize = 8'd39;
        8'd132: linearize = 8'd40;
        8'd133: linearize = 8'd41;
        8'd134: linearize = 8'd42;
        8'd135: linearize = 8'd43;
        8'd136: linearize = 8'd44;
        8'd137: linearize = 8'd45;
        8'd138: linearize = 8'd46;
        8'd139: linearize = 8'd47;
        8'd140: linearize = 8'd48;
        8'd141: linearize = 8'd49;
        8'd142: linearize = 8'd50;
        8'd143: linearize = 8'd50;
        8'd144: linearize = 8'd51;
        8'd145: linearize = 8'd52;
        8'd146: linearize = 8'd54;
        8'd147: linearize = 8'd55;
        8'd148: linearize = 8'd56;
        8'd149: linearize = 8'd57;
        8'd150: linearize = 8'd58;
        8'd151: linearize = 8'd59;
        8'd152: linearize = 8'd60;
        8'd153: linearize = 8'd61;
        8'd154: linearize = 8'd62;
        8'd155: linearize = 8'd63;
        8'd156: linearize = 8'd64;
        8'd157: linearize = 8'd66;
        8'd158: linearize = 8'd67;
        8'd159: linearize = 8'd68;
        8'd160: linearize = 8'd69;
        8'd161: linearize = 8'd70;
        8'd162: linearize = 8'd72;
        8'd163: linearize = 8'd73;
        8'd164: linearize = 8'd74;
        8'd165: linearize = 8'd75;
        8'd166: linearize = 8'd77;
        8'd167: linearize = 8'd78;
        8'd168: linearize = 8'd79;
        8'd169: linearize = 8'd81;
        8'd170: linearize = 8'd82;
        8'd171: linearize = 8'd83;
        8'd172: linearize = 8'd85;
        8'd173: linearize = 8'd86;
        8'd174: linearize = 8'd87;
        8'd175: linearize = 8'd89;
        8'd176: linearize = 8'd90;
        8'd177: linearize = 8'd92;
        8'd178: linearize = 8'd93;
        8'd179: linearize = 8'd95;
        8'd180: linearize = 8'd96;
        8'd181: linearize = 8'd98;
        8'd182: linearize = 8'd99;
        8'd183: linearize = 8'd101;
        8'd184: linearize = 8'd102;
        8'd185: linearize = 8'd104;
        8'd186: linearize = 8'd105;
        8'd187: linearize = 8'd107;
        8'd188: linearize = 8'd109;
        8'd189: linearize = 8'd110;
        8'd190: linearize = 8'd112;
        8'd191: linearize = 8'd114;
        8'd192: linearize = 8'd115;
        8'd193: linearize = 8'd117;
        8'd194: linearize = 8'd119;
        8'd195: linearize = 8'd120;
        8'd196: linearize = 8'd122;
        8'd197: linearize = 8'd124;
        8'd198: linearize = 8'd126;
        8'd199: linearize = 8'd127;
        8'd200: linearize = 8'd129;
        8'd201: linearize = 8'd131;
        8'd202: linearize = 8'd133;
        8'd203: linearize = 8'd135;
        8'd204: linearize = 8'd137;
        8'd205: linearize = 8'd138;
        8'd206: linearize = 8'd140;
        8'd207: linearize = 8'd142;
        8'd208: linearize = 8'd144;
        8'd209: linearize = 8'd146;
        8'd210: linearize = 8'd148;
        8'd211: linearize = 8'd150;
        8'd212: linearize = 8'd152;
        8'd213: linearize = 8'd154;
        8'd214: linearize = 8'd156;
        8'd215: linearize = 8'd158;
        8'd216: linearize = 8'd160;
        8'd217: linearize = 8'd162;
        8'd218: linearize = 8'd164;
        8'd219: linearize = 8'd167;
        8'd220: linearize = 8'd169;
        8'd221: linearize = 8'd171;
        8'd222: linearize = 8'd173;
        8'd223: linearize = 8'd175;
        8'd224: linearize = 8'd177;
        8'd225: linearize = 8'd180;
        8'd226: linearize = 8'd182;
        8'd227: linearize = 8'd184;
        8'd228: linearize = 8'd186;
        8'd229: linearize = 8'd189;
        8'd230: linearize = 8'd191;
        8'd231: linearize = 8'd193;
        8'd232: linearize = 8'd196;
        8'd233: linearize = 8'd198;
        8'd234: linearize = 8'd200;
        8'd235: linearize = 8'd203;
        8'd236: linearize = 8'd205;
        8'd237: linearize = 8'd208;
        8'd238: linearize = 8'd210;
        8'd239: linearize = 8'd213;
        8'd240: linearize = 8'd215;
        8'd241: linearize = 8'd218;
        8'd242: linearize = 8'd220;
        8'd243: linearize = 8'd223;
        8'd244: linearize = 8'd225;
        8'd245: linearize = 8'd228;
        8'd246: linearize = 8'd231;
        8'd247: linearize = 8'd233;
        8'd248: linearize = 8'd236;
        8'd249: linearize = 8'd239;
        8'd250: linearize = 8'd241;
        8'd251: linearize = 8'd244;
        8'd252: linearize = 8'd247;
        8'd253: linearize = 8'd249;
        8'd254: linearize = 8'd252;
        8'd255: linearize = 8'd255;
    endcase
endfunction

`endif
